//SystemVerilog
module rom_pipelined #(parameter STAGES=2)(
    input clk,
    input [9:0] addr_in,
    output [7:0] data_out
);
    reg [9:0] pipe_addr [0:STAGES-1];
    reg [7:0] pipe_data [0:STAGES-1];
    reg [7:0] mem [0:1023];
    
    integer i;
    
    // Initialize memory with some default values
    initial begin
        for (i = 0; i < 1024; i = i + 1)
            mem[i] = i & 8'hFF; // Simple pattern for testing
    end
    
    always @(posedge clk) begin
        // Move the first register for addr_in after the combinational logic
        pipe_data[0] <= mem[addr_in]; // Directly use addr_in for data retrieval
        for(i = 1; i < STAGES; i = i + 1)
            pipe_data[i] <= pipe_data[i-1];

        // Update pipe_addr after data processing
        pipe_addr[0] <= addr_in; // Keep the addr_in register
        for(i = 1; i < STAGES; i = i + 1)
            pipe_addr[i] <= pipe_addr[i-1];
    end
    
    assign data_out = pipe_data[STAGES-1];
endmodule