module Adder_1(
    input [3:0] A,
    input [3:0] B,
    output [4:0] sum
);
    assign sum = A + B;
endmodule