module dual_hamming_encoder(
    input clk, rst_n,
    input [3:0] data_a, data_b,
    output reg [6:0] encoded_a, encoded_b
);
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            encoded_a <= 7'b0;
            encoded_b <= 7'b0;
        end else begin
            // Channel A
            encoded_a[0] <= data_a[0] ^ data_a[1] ^ data_a[3];
            encoded_a[1] <= data_a[0] ^ data_a[2] ^ data_a[3];
            encoded_a[2] <= data_a[0];
            encoded_a[3] <= data_a[1] ^ data_a[2] ^ data_a[3];
            encoded_a[4] <= data_a[1];
            encoded_a[5] <= data_a[2];
            encoded_a[6] <= data_a[3];
            
            // Channel B
            encoded_b[0] <= data_b[0] ^ data_b[1] ^ data_b[3];
            encoded_b[1] <= data_b[0] ^ data_b[2] ^ data_b[3];
            encoded_b[2] <= data_b[0];
            encoded_b[3] <= data_b[1] ^ data_b[2] ^ data_b[3];
            encoded_b[4] <= data_b[1];
            encoded_b[5] <= data_b[2];
            encoded_b[6] <= data_b[3];
        end
    end
endmodule