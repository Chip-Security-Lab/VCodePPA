module nand_xor_gate (
    input wire A, B, C,   // 输入A, B, C
    output wire Y         // 输出Y
);
    assign Y = ~(A & B) ^ C;
endmodule
