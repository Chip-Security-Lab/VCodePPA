//SystemVerilog
// Submodule to generate Propagate (P) and Generate (G) signals
module pg_generator (
    input [3:0] a,
    input [3:0] b,
    output [3:0] p, // Pi = Ai XOR Bi
    output [3:0] g  // Gi = Ai AND Bi
);

  genvar i;
  generate
    for (i = 0; i < 4; i = i + 1) begin : gen_pg_logic
      assign p[i] = a[i] ^ b[i];
      assign g[i] = a[i] & b[i];
    end
  endgenerate

endmodule

// Submodule for Carry Lookahead Logic
module carry_lookahead (
    input [3:0] p, // Propagate signals
    input [3:0] g, // Generate signals
    input       cin,
    output [4:0] c  // Carry signals: c[0] is cin, c[i+1] is carry into bit i, c[4] is cout
);

  assign c[0] = cin;
  assign c[1] = g[0] | (p[0] & c[0]);
  assign c[2] = g[1] | (p[1] & g[0]) | (p[1] & p[0] & c[0]);
  assign c[3] = g[2] | (p[2] & g[1]) | (p[2] & p[1] & g[0]) | (p[2] & p[1] & p[0] & c[0]);
  assign c[4] = g[3] | (p[3] & g[2]) | (p[3] & p[2] & g[1]) | (p[3] & p[2] & p[1] & g[0]) | (p[3] & p[2] & p[1] & p[0] & c[0]);

endmodule

// Submodule to generate Sum signals
module sum_generator (
    input [3:0] p, // Propagate signals
    input [3:0] c, // Carry signals (c[0] to c[3])
    output [3:0] sum // Sum signals: Sum[i] = Pi XOR C[i]
);

  genvar i;
  generate
    for (i = 0; i < 4; i = i + 1) begin : gen_sum_logic
      assign sum[i] = p[i] ^ c[i];
    end
  endgenerate

endmodule

// Refactored 4-bit Carry-Lookahead Adder (CLA) block using submodules
module cla_4bit (
    input [3:0] a,
    input [3:0] b,
    input       cin,
    output [3:0] sum,
    output      cout // Carry out of bit 3
);

  wire [3:0] p; // Propagate signals
  wire [3:0] g; // Generate signals
  wire [4:0] c; // Carry signals (c[0] is cin, c[4] is cout)

  // Instantiate PG generator submodule
  pg_generator u_pg_gen (
      .a(a),
      .b(b),
      .p(p),
      .g(g)
  );

  // Instantiate Carry Lookahead submodule
  carry_lookahead u_cla_logic (
      .p(p),
      .g(g),
      .cin(cin),
      .c(c)
  );

  // Instantiate Sum generator submodule
  sum_generator u_sum_gen (
      .p(p),
      .c(c[3:0]), // Connect relevant carries (c[0] to c[3])
      .sum(sum)
  );

  // Output carry is the last carry generated by the CLA logic
  assign cout = c[4];

endmodule


// Top-level 8-bit adder module using hierarchical 4-bit CLA blocks
// Original module name retained, ports updated for 8-bit operation with carry
module adder_2 (
    input [7:0] a,
    input [7:0] b,
    input       cin,
    output [7:0] sum,
    output      cout
);

  wire c4; // Carry out of the lower 4 bits (bit 3), carry into the upper 4 bits (bit 4)

  // Instantiate the lower 4-bit CLA block (bits 3 down to 0)
  cla_4bit u_cla_low (
      .a   (a[3:0]),
      .b   (b[3:0]),
      .cin (cin),
      .sum (sum[3:0]),
      .cout(c4)
  );

  // Instantiate the upper 4-bit CLA block (bits 7 down to 4)
  cla_4bit u_cla_high (
      .a   (a[7:4]),
      .b   (b[7:4]),
      .cin (c4), // Connect carry-out of lower block to carry-in of upper block
      .sum (sum[7:4]),
      .cout(cout) // Carry-out of upper block is the final cout
  );

endmodule