//SystemVerilog
module ParityLatch #(parameter DW=7) (
    input clk, en,
    input [DW-1:0] data,
    output reg [DW:0] q
);

// LUT-based parity calculation
reg [DW:0] lut_parity [0:255];

initial begin
    lut_parity[0] = 0;
    lut_parity[1] = 1;
    lut_parity[2] = 1;
    lut_parity[3] = 0;
    lut_parity[4] = 1;
    lut_parity[5] = 0;
    lut_parity[6] = 0;
    lut_parity[7] = 1;
    lut_parity[8] = 1;
    lut_parity[9] = 0;
    lut_parity[10] = 0;
    lut_parity[11] = 1;
    lut_parity[12] = 0;
    lut_parity[13] = 1;
    lut_parity[14] = 1;
    lut_parity[15] = 0;
    lut_parity[16] = 1;
    lut_parity[17] = 0;
    lut_parity[18] = 0;
    lut_parity[19] = 1;
    lut_parity[20] = 0;
    lut_parity[21] = 1;
    lut_parity[22] = 1;
    lut_parity[23] = 0;
    lut_parity[24] = 0;
    lut_parity[25] = 1;
    lut_parity[26] = 1;
    lut_parity[27] = 0;
    lut_parity[28] = 1;
    lut_parity[29] = 0;
    lut_parity[30] = 0;
    lut_parity[31] = 1;
    lut_parity[32] = 1;
    lut_parity[33] = 0;
    lut_parity[34] = 0;
    lut_parity[35] = 1;
    lut_parity[36] = 0;
    lut_parity[37] = 1;
    lut_parity[38] = 1;
    lut_parity[39] = 0;
    lut_parity[40] = 0;
    lut_parity[41] = 1;
    lut_parity[42] = 1;
    lut_parity[43] = 0;
    lut_parity[44] = 1;
    lut_parity[45] = 0;
    lut_parity[46] = 0;
    lut_parity[47] = 1;
    lut_parity[48] = 0;
    lut_parity[49] = 1;
    lut_parity[50] = 1;
    lut_parity[51] = 0;
    lut_parity[52] = 1;
    lut_parity[53] = 0;
    lut_parity[54] = 0;
    lut_parity[55] = 1;
    lut_parity[56] = 1;
    lut_parity[57] = 0;
    lut_parity[58] = 0;
    lut_parity[59] = 1;
    lut_parity[60] = 0;
    lut_parity[61] = 1;
    lut_parity[62] = 1;
    lut_parity[63] = 0;
    lut_parity[64] = 1;
    lut_parity[65] = 0;
    lut_parity[66] = 0;
    lut_parity[67] = 1;
    lut_parity[68] = 0;
    lut_parity[69] = 1;
    lut_parity[70] = 1;
    lut_parity[71] = 0;
    lut_parity[72] = 0;
    lut_parity[73] = 1;
    lut_parity[74] = 1;
    lut_parity[75] = 0;
    lut_parity[76] = 1;
    lut_parity[77] = 0;
    lut_parity[78] = 0;
    lut_parity[79] = 1;
    lut_parity[80] = 0;
    lut_parity[81] = 1;
    lut_parity[82] = 1;
    lut_parity[83] = 0;
    lut_parity[84] = 1;
    lut_parity[85] = 0;
    lut_parity[86] = 0;
    lut_parity[87] = 1;
    lut_parity[88] = 1;
    lut_parity[89] = 0;
    lut_parity[90] = 0;
    lut_parity[91] = 1;
    lut_parity[92] = 0;
    lut_parity[93] = 1;
    lut_parity[94] = 1;
    lut_parity[95] = 0;
    lut_parity[96] = 0;
    lut_parity[97] = 1;
    lut_parity[98] = 1;
    lut_parity[99] = 0;
    lut_parity[100] = 1;
    lut_parity[101] = 0;
    lut_parity[102] = 0;
    lut_parity[103] = 1;
    lut_parity[104] = 1;
    lut_parity[105] = 0;
    lut_parity[106] = 0;
    lut_parity[107] = 1;
    lut_parity[108] = 0;
    lut_parity[109] = 1;
    lut_parity[110] = 1;
    lut_parity[111] = 0;
    lut_parity[112] = 1;
    lut_parity[113] = 0;
    lut_parity[114] = 0;
    lut_parity[115] = 1;
    lut_parity[116] = 0;
    lut_parity[117] = 1;
    lut_parity[118] = 1;
    lut_parity[119] = 0;
    lut_parity[120] = 0;
    lut_parity[121] = 1;
    lut_parity[122] = 1;
    lut_parity[123] = 0;
    lut_parity[124] = 1;
    lut_parity[125] = 0;
    lut_parity[126] = 0;
    lut_parity[127] = 1;
    lut_parity[128] = 1;
    lut_parity[129] = 0;
    lut_parity[130] = 0;
    lut_parity[131] = 1;
    lut_parity[132] = 0;
    lut_parity[133] = 1;
    lut_parity[134] = 1;
    lut_parity[135] = 0;
    lut_parity[136] = 0;
    lut_parity[137] = 1;
    lut_parity[138] = 1;
    lut_parity[139] = 0;
    lut_parity[140] = 1;
    lut_parity[141] = 0;
    lut_parity[142] = 0;
    lut_parity[143] = 1;
    lut_parity[144] = 0;
    lut_parity[145] = 1;
    lut_parity[146] = 1;
    lut_parity[147] = 0;
    lut_parity[148] = 1;
    lut_parity[149] = 0;
    lut_parity[150] = 0;
    lut_parity[151] = 1;
    lut_parity[152] = 1;
    lut_parity[153] = 0;
    lut_parity[154] = 0;
    lut_parity[155] = 1;
    lut_parity[156] = 0;
    lut_parity[157] = 1;
    lut_parity[158] = 1;
    lut_parity[159] = 0;
    lut_parity[160] = 0;
    lut_parity[161] = 1;
    lut_parity[162] = 1;
    lut_parity[163] = 0;
    lut_parity[164] = 1;
    lut_parity[165] = 0;
    lut_parity[166] = 0;
    lut_parity[167] = 1;
    lut_parity[168] = 1;
    lut_parity[169] = 0;
    lut_parity[170] = 0;
    lut_parity[171] = 1;
    lut_parity[172] = 0;
    lut_parity[173] = 1;
    lut_parity[174] = 1;
    lut_parity[175] = 0;
    lut_parity[176] = 0;
    lut_parity[177] = 1;
    lut_parity[178] = 1;
    lut_parity[179] = 0;
    lut_parity[180] = 1;
    lut_parity[181] = 0;
    lut_parity[182] = 0;
    lut_parity[183] = 1;
    lut_parity[184] = 1;
    lut_parity[185] = 0;
    lut_parity[186] = 0;
    lut_parity[187] = 1;
    lut_parity[188] = 0;
    lut_parity[189] = 1;
    lut_parity[190] = 1;
    lut_parity[191] = 0;
    lut_parity[192] = 0;
    lut_parity[193] = 1;
    lut_parity[194] = 1;
    lut_parity[195] = 0;
    lut_parity[196] = 1;
    lut_parity[197] = 0;
    lut_parity[198] = 0;
    lut_parity[199] = 1;
    lut_parity[200] = 1;
    lut_parity[201] = 0;
    lut_parity[202] = 0;
    lut_parity[203] = 1;
    lut_parity[204] = 0;
    lut_parity[205] = 1;
    lut_parity[206] = 1;
    lut_parity[207] = 0;
    lut_parity[208] = 0;
    lut_parity[209] = 1;
    lut_parity[210] = 1;
    lut_parity[211] = 0;
    lut_parity[212] = 1;
    lut_parity[213] = 0;
    lut_parity[214] = 0;
    lut_parity[215] = 1;
    lut_parity[216] = 1;
    lut_parity[217] = 0;
    lut_parity[218] = 0;
    lut_parity[219] = 1;
    lut_parity[220] = 0;
    lut_parity[221] = 1;
    lut_parity[222] = 1;
    lut_parity[223] = 0;
    lut_parity[224] = 0;
    lut_parity[225] = 1;
    lut_parity[226] = 1;
    lut_parity[227] = 0;
    lut_parity[228] = 1;
    lut_parity[229] = 0;
    lut_parity[230] = 0;
    lut_parity[231] = 1;
    lut_parity[232] = 1;
    lut_parity[233] = 0;
    lut_parity[234] = 0;
    lut_parity[235] = 1;
    lut_parity[236] = 0;
    lut_parity[237] = 1;
    lut_parity[238] = 1;
    lut_parity[239] = 0;
    lut_parity[240] = 0;
    lut_parity[241] = 1;
    lut_parity[242] = 1;
    lut_parity[243] = 0;
    lut_parity[244] = 1;
    lut_parity[245] = 0;
    lut_parity[246] = 0;
    lut_parity[247] = 1;
    lut_parity[248] = 1;
    lut_parity[249] = 0;
    lut_parity[250] = 0;
    lut_parity[251] = 1;
    lut_parity[252] = 0;
    lut_parity[253] = 1;
    lut_parity[254] = 1;
    lut_parity[255] = 0;
end

always @(posedge clk)
    if(en) q <= {lut_parity[data], data};

endmodule