module adder_7 (a, b, sum);
  input a, b;
  output sum;
  assign sum = a + b;
endmodule