//SystemVerilog
// SystemVerilog
module rr_async_icmu (
    input rst,
    input [7:0] interrupt_in,
    input ctx_save_done,
    output reg [7:0] int_grant,
    output reg [2:0] int_vector,
    output reg context_save_req
);
    reg [2:0] last_served;
    reg [7:0] masked_ints;

    // Reorganized combinatorial logic
    always @(*) begin
        masked_ints = interrupt_in;
        context_save_req = |masked_ints;

        // Use function call
        int_grant = select_next(masked_ints, last_served);
        int_vector = encode_vec(int_grant);
    end

    always @(posedge ctx_save_done or posedge rst) begin
        if (rst) begin
            last_served <= 3'b0;
        end else begin
            last_served <= int_vector;
        end
    end

    // 3-bit borrow-based subtractor function
    // Computes a - b, returns {BorrowOut, Difference}
    function automatic [3:0] subtractor_3bit;
        input [2:0] a;
        input [2:0] b;
        reg [2:0] diff;
        reg [2:0] bout_chain; // Internal borrow chain

        begin
            // Bit 0 (LSB)
            diff[0] = a[0] ^ b[0] ^ 1'b0; // Assume Bin = 0 for A - B
            bout_chain[0] = (~a[0] & b[0]) | (~a[0] & 1'b0) | (b[0] & 1'b0);

            // Bit 1
            diff[1] = a[1] ^ b[1] ^ bout_chain[0];
            bout_chain[1] = (~a[1] & b[1]) | (~a[1] & bout_chain[0]) | (b[1] & bout_chain[0]);

            // Bit 2 (MSB)
            diff[2] = a[2] ^ b[2] ^ bout_chain[1];
            bout_chain[2] = (~a[2] & b[2]) | (~a[2] & bout_chain[1]) | (b[2] & bout_chain[1]);

            // BorrowOut is the borrow generated by the MSB stage
            subtractor_3bit = {bout_chain[2], diff};
        end
    endfunction


    // Modified function implementation with borrow-based subtractor for mask
    function [7:0] select_next;
        input [7:0] ints;
        input [2:0] last;
        reg [7:0] mask, high_result, any_result;
        integer i;
        reg [2:0] i_3bit;
        reg [3:0] sub_result; // {BorrowOut, Diff}
        reg borrow_out;

        begin
            mask = 0;
            high_result = 0;
            any_result = 0;

            // Create mask using borrow-based subtractor for comparison (i > last)
            // i > last is equivalent to last < i
            // last < i is equivalent to borrow_out of (last - i) being 1
            for (i = 0; i < 8; i = i + 1) begin
                i_3bit = i; // Cast integer i to 3 bits

                // Compute last - i_3bit using borrow-based subtractor
                sub_result = subtractor_3bit(last, i_3bit);
                borrow_out = sub_result[3]; // BorrowOut is the MSB

                if (borrow_out) begin // If last < i_3bit (i.e., i > last)
                    mask[i] = 1'b1;
                end else begin
                    mask[i] = 1'b0;
                end
            end

            // Find interrupts higher than last using mask
            high_result = ints & mask;

            // Find all interrupts
            any_result = ints;

            // Select result (already in this format)
            if (|high_result) begin
                select_next = high_result;
            end else begin
                select_next = any_result;
            end
        end
    endfunction

    function [2:0] encode_vec;
        input [7:0] grant;
        begin
            casez(grant)
                8'b???????1: encode_vec = 3'd0;
                8'b??????10: encode_vec = 3'd1;
                8'b?????100: encode_vec = 3'd2;
                8'b????1000: encode_vec = 3'd3;
                8'b???10000: encode_vec = 3'd4;
                8'b??100000: encode_vec = 3'd5;
                8'b?1000000: encode_vec = 3'd6;
                8'b10000000: encode_vec = 3'd7;
                default: encode_vec = 3'd0;
            endcase
        end
    endfunction

    function [2:0] find_first;
        input [7:0] val;
        begin
            casez(val)
                8'b???????1: find_first = 3'd0;
                8'b??????10: find_first = 3'd1;
                8'b?????100: find_first = 3'd2;
                8'b????1000: find_first = 3'd3;
                8'b???10000: find_first = 3'd4;
                8'b??100000: find_first = 3'd5;
                8'b?1000000: find_first = 3'd6;
                8'b10000000: find_first = 3'd7;
                default: find_first = 3'd0;
            endcase
        end
    endfunction
endmodule