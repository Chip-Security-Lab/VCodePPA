module LevelITRC #(parameter CHANNELS=4, TIMEOUT=8) (
    input clk, rst,
    input [CHANNELS-1:0] level_irq,
    output reg irq_valid,
    output reg [$clog2(CHANNELS)-1:0] active_channel
);
    reg [CHANNELS-1:0] irq_active;
    reg [$clog2(TIMEOUT):0] timeout_counter [0:CHANNELS-1];
    integer i;
    
    always @(posedge clk) begin
        if (rst) begin
            irq_active <= 0;
            irq_valid <= 0;
            active_channel <= 0;
            for (i = 0; i < CHANNELS; i = i + 1)
                timeout_counter[i] <= 0;
        end else begin
            // Process each channel individually
            if (level_irq[0] && !irq_active[0]) begin
                irq_active[0] <= 1;
                timeout_counter[0] <= TIMEOUT;
            end else if (irq_active[0] && timeout_counter[0] > 0) begin
                timeout_counter[0] <= timeout_counter[0] - 1;
            end else if (irq_active[0]) begin
                irq_active[0] <= 0; // Auto-clear after timeout
            end
            
            if (level_irq[1] && !irq_active[1]) begin
                irq_active[1] <= 1;
                timeout_counter[1] <= TIMEOUT;
            end else if (irq_active[1] && timeout_counter[1] > 0) begin
                timeout_counter[1] <= timeout_counter[1] - 1;
            end else if (irq_active[1]) begin
                irq_active[1] <= 0;
            end
            
            if (level_irq[2] && !irq_active[2]) begin
                irq_active[2] <= 1;
                timeout_counter[2] <= TIMEOUT;
            end else if (irq_active[2] && timeout_counter[2] > 0) begin
                timeout_counter[2] <= timeout_counter[2] - 1;
            end else if (irq_active[2]) begin
                irq_active[2] <= 0;
            end
            
            if (level_irq[3] && !irq_active[3]) begin
                irq_active[3] <= 1;
                timeout_counter[3] <= TIMEOUT;
            end else if (irq_active[3] && timeout_counter[3] > 0) begin
                timeout_counter[3] <= timeout_counter[3] - 1;
            end else if (irq_active[3]) begin
                irq_active[3] <= 0;
            end
            
            // Find highest priority active interrupt
            irq_valid <= |irq_active;
            if (irq_active[3]) active_channel <= 2'd3;
            else if (irq_active[2]) active_channel <= 2'd2;
            else if (irq_active[1]) active_channel <= 2'd1;
            else if (irq_active[0]) active_channel <= 2'd0;
        end
    end
endmodule