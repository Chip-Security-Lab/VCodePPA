module or_gate_2input_1bit (
    input wire a,
    input wire b,
    output wire y
);
    assign y = a | b;
endmodule
