module xor_alias(
    input in1, 
    input in2,
    output result
);
    assign result = in1 ^ in2;
endmodule