// 单行注释
module adder_5 (input a, b, output sum);
    // Assign statement
    assign sum = a + b;
    // End of module
endmodule