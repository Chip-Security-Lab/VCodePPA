module not_gate_1bit (
    input wire A,
    output wire Y
);
    assign Y = ~A;
endmodule
