module adder_12 (input a, b, output sum);
  // This is an example of a basic adder
  assign sum = a + b; // Main add operation
endmodule