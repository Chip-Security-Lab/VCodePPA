//SystemVerilog
// IEEE 1364-2005 Verilog标准
module prio_enc_function #(parameter W=16)(
  input [W-1:0] req,
  output reg [$clog2(W)-1:0] enc_addr
);

  // 使用组合逻辑查找最高优先级位置
  always @(*) begin
    enc_addr = 0;
    casez(req)
      16'b1???????????????: enc_addr = 4'd15;
      16'b01??????????????: enc_addr = 4'd14;
      16'b001?????????????: enc_addr = 4'd13;
      16'b0001????????????: enc_addr = 4'd12;
      16'b00001???????????: enc_addr = 4'd11;
      16'b000001??????????: enc_addr = 4'd10;
      16'b0000001?????????: enc_addr = 4'd9;
      16'b00000001????????: enc_addr = 4'd8;
      16'b000000001???????: enc_addr = 4'd7;
      16'b0000000001??????: enc_addr = 4'd6;
      16'b00000000001?????: enc_addr = 4'd5;
      16'b000000000001????: enc_addr = 4'd4;
      16'b0000000000001???: enc_addr = 4'd3;
      16'b00000000000001??: enc_addr = 4'd2;
      16'b000000000000001?: enc_addr = 4'd1;
      16'b0000000000000001: enc_addr = 4'd0;
      default:              enc_addr = 4'd0;
    endcase
  end

endmodule