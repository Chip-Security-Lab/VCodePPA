module OR_basic(
    input a, b,
    output y
);
    assign y = a | b;  // 基本逻辑或操作
endmodule
