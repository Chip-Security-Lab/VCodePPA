module Triple_AND(
    input a, b, c,
    output out
);
    assign out = a & b & c; // 三输入逻辑与
endmodule
