module adder_1 (input a, b, output sum);
  assign sum = a + b;
endmodule