module xor2_1 (
    input wire A, B,
    output wire Y
);
    assign Y = A ^ B; // 基本的2输入异或门
endmodule
