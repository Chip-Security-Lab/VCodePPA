module moore_3state_mem_write_ctrl #(parameter ADDR_WIDTH = 4)(
  input  clk,
  input  rst,
  input  start,
  output reg we,
  output reg [ADDR_WIDTH-1:0] addr
);
  reg [1:0] state, next_state;
  localparam IDLE    = 2'b00,
             SET_ADDR= 2'b01,
             WRITE   = 2'b10;

  always @(posedge clk or posedge rst) begin
    if (rst) begin
      state <= IDLE;
      addr  <= 0;
    end else begin
      state <= next_state;
      if (state == SET_ADDR) addr <= addr + 1;
    end
  end

  always @* begin
    we = 1'b0;
    case (state)
      IDLE:    next_state = start ? SET_ADDR : IDLE;
      SET_ADDR:next_state = WRITE;
      WRITE:   next_state = IDLE;
    endcase
    // Moore输出：只有在当前状态为WRITE时才置we=1
    if (state == WRITE) we = 1'b1;
  end
endmodule
