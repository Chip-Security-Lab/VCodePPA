/*
 * Multi-line comment
 * This is a simple adder module
 */
module adder_6 (input a, b, output sum);
  assign sum = a + b;
endmodule