module adder_3 (input wire a, input wire b, output wire sum);
  assign sum = a + b;
endmodule