//SystemVerilog
module pipeline_arbiter(
  input wire clk, async_reset_n,
  input wire [3:0] request,
  input wire ready,
  output reg [3:0] grant,
  output reg valid
);
  reg [3:0] req_stage1, req_stage2;
  reg [1:0] state, next_state;
  reg valid_pending;
  
  always @(posedge clk or negedge async_reset_n) begin
    if (!async_reset_n) begin
      state <= 2'b00; 
      req_stage1 <= 4'b0; 
      req_stage2 <= 4'b0; 
      grant <= 4'b0; 
      valid <= 1'b0;
      valid_pending <= 1'b0;
    end else begin
      state <= next_state;
      req_stage1 <= request;
      req_stage2 <= req_stage1;
      
      if (valid_pending && ready) begin
        valid_pending <= 1'b0;
        valid <= 1'b0;
      end else if (|request && !valid_pending) begin
        valid_pending <= 1'b1;
        valid <= 1'b1;
      end
      
      // Pipelined arbitration logic
    end
  end
endmodule