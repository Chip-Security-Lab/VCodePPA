//SystemVerilog
module MedianFilter #(parameter WIDTH=8) (
    input [WIDTH-1:0] a, b, c,
    output reg [WIDTH-1:0] med
);
    reg [WIDTH-1:0] max_ab;
    reg [WIDTH-1:0] min_ab;
    reg [1:0] comp_result;
    
    always @(*) begin
        // 使用比较结果位表示a与b的关系
        comp_result[0] = (a > b);  // a是否大于b
        comp_result[1] = (a < b);  // a是否小于b
        
        // 使用case语句确定max_ab和min_ab
        case(comp_result)
            2'b01: begin  // a < b
                max_ab = b;
                min_ab = a;
            end
            2'b10: begin  // a > b
                max_ab = a;
                min_ab = b;
            end
            default: begin  // a == b
                max_ab = a;
                min_ab = a;
            end
        endcase
        
        // 使用case语句确定中值
        casez({c > max_ab, c < min_ab})
            2'b1?: med = max_ab;  // c > max_ab
            2'b01: med = min_ab;  // c < min_ab
            default: med = c;     // min_ab <= c <= max_ab
        endcase
    end
endmodule