module not_gate_comb (
    input wire A,
    output wire Y
);
    assign Y = ~A;
endmodule
