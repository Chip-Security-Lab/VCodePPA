module async_mult (
    input [3:0] A, B,
    output [7:0] P,
    input start,
    output done
);
    // 异步状态机实现
    reg [2:0] state;
    reg [3:0] multiplicand;
    reg [3:0] multiplier;
    reg [7:0] product;
    reg done_reg;
    
    parameter IDLE = 3'b000;
    parameter INIT = 3'b001;
    parameter ADD = 3'b010;
    parameter SHIFT = 3'b011;
    parameter FINISH = 3'b100;
    
    reg [2:0] counter;
    
    // 状态转换逻辑
    always @(state or start or counter or multiplier[0]) begin
        case(state)
            IDLE: state = start ? INIT : IDLE;
            INIT: state = ADD;
            ADD: state = SHIFT;
            SHIFT: state = (counter == 3'b011) ? FINISH : ADD;
            FINISH: state = IDLE;
            default: state = IDLE;
        endcase
    end
    
    // 数据处理逻辑
    always @(state) begin
        case(state)
            IDLE: begin
                done_reg = 1'b1;
                counter = 3'b000;
            end
            
            INIT: begin
                multiplicand = A;
                multiplier = B;
                product = 8'b0;
                counter = 3'b000;
                done_reg = 1'b0;
            end
            
            ADD: begin
                if(multiplier[0])
                    product[7:4] = product[7:4] + multiplicand;
            end
            
            SHIFT: begin
                multiplier = multiplier >> 1;
                product = product >> 1;
                counter = counter + 1;
            end
            
            FINISH: begin
                done_reg = 1'b1;
            end
        endcase
    end
    
    assign P = product;
    assign done = done_reg;
endmodule