//SystemVerilog
module pwm_div #(parameter HIGH=3, LOW=5) (
    input clk, rst_n,
    output reg out
);
    reg [7:0] cnt;
    reg cnt_is_high;
    
    always @(posedge clk) begin
        if(!rst_n) begin
            cnt <= 0;
            cnt_is_high <= 0;
        end else begin
            cnt <= (cnt == HIGH+LOW-1) ? 0 : cnt + 1;
            cnt_is_high <= (cnt + 1 < HIGH) || ((cnt == HIGH+LOW-1) && (HIGH > 0));
        end
    end
    
    always @(posedge clk) begin
        if(!rst_n) begin
            out <= 0;
        end else begin
            out <= cnt_is_high;
        end
    end
endmodule