//SystemVerilog
module usb_isoc_manager #(
    parameter NUM_ENDPOINTS = 4,
    parameter DATA_WIDTH = 16
)(
    input wire clock, reset_b,
    input wire sof_received,
    input wire [10:0] frame_number,
    input wire [3:0] endpoint_select,
    input wire transfer_ready,
    input wire [DATA_WIDTH-1:0] tx_data,
    output reg transfer_active,
    output reg [DATA_WIDTH-1:0] rx_data,
    output reg [NUM_ENDPOINTS-1:0] endpoint_status,
    output reg [1:0] bandwidth_state
);
    // Bandwidth reservation states
    localparam IDLE = 2'b00;
    localparam RESERVED = 2'b01;
    localparam ACTIVE = 2'b10;
    localparam COMPLETE = 2'b11;
    
    // Per-endpoint configuration and state
    reg [2:0] interval [0:NUM_ENDPOINTS-1];
    reg [10:0] last_frame [0:NUM_ENDPOINTS-1];
    reg [10:0] frame_diff [0:NUM_ENDPOINTS-1]; // Precompute frame differences
    
    integer i;
    always @(posedge clock or negedge reset_b) begin
        if (!reset_b) begin
            transfer_active <= 1'b0;
            bandwidth_state <= IDLE;
            endpoint_status <= {NUM_ENDPOINTS{1'b0}};
            for (i = 0; i < NUM_ENDPOINTS; i = i + 1) begin
                interval[i] <= 3'd1;         // Default interval of 1 frame
                last_frame[i] <= 11'h7FF;    // Invalid frame number
                frame_diff[i] <= 11'd0;      // Initialize difference
            end
        end else if (sof_received) begin
            // Precompute all frame differences in parallel
            for (i = 0; i < NUM_ENDPOINTS; i = i + 1) begin
                frame_diff[i] <= frame_number - last_frame[i];
            end
            
            // Use the precomputed differences for comparison
            for (i = 0; i < NUM_ENDPOINTS; i = i + 1) begin
                // Simplify comparison by checking only relevant bits
                // and avoid unnecessary zero-extension
                endpoint_status[i] <= (frame_diff[i][2:0] >= interval[i]);
            end
        end
    end
endmodule