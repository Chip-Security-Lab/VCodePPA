module Sub1(input [7:0] a,b, output [7:0] result);
    assign result = a - b;
endmodule