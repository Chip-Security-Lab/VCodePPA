module eth_checksum_verifier (
    input wire clock,
    input wire reset,
    input wire data_valid,
    input wire [7:0] rx_byte,
    input wire packet_start,
    input wire packet_end,
    output reg checksum_ok,
    output reg checksum_valid
);
    reg [15:0] checksum;
    reg [15:0] computed_checksum;
    reg [2:0] state;
    reg [9:0] byte_count;
    
    localparam IDLE = 3'd0, HEADER = 3'd1, DATA = 3'd2, CHECKSUM_L = 3'd3, CHECKSUM_H = 3'd4;
    
    always @(posedge clock or posedge reset) begin
        if (reset) begin
            state <= IDLE;
            byte_count <= 10'd0;
            checksum <= 16'd0;
            computed_checksum <= 16'd0;
            checksum_ok <= 1'b0;
            checksum_valid <= 1'b0;
        end else begin
            if (packet_start) begin
                state <= HEADER;
                byte_count <= 10'd0;
                computed_checksum <= 16'd0;
                checksum_ok <= 1'b0;
                checksum_valid <= 1'b0;
            end else if (data_valid) begin
                case (state)
                    HEADER: begin
                        if (byte_count < 13) begin
                            byte_count <= byte_count + 1'b1;
                        end else begin
                            state <= DATA;
                            byte_count <= 10'd0;
                        end
                    end
                    
                    DATA: begin
                        // Sum all data bytes for simple checksum calculation
                        computed_checksum <= computed_checksum + rx_byte;
                        
                        // Assume checksum is last 2 bytes of packet
                        if (packet_end) begin
                            state <= CHECKSUM_L;
                        end
                    end
                    
                    CHECKSUM_L: begin
                        checksum[7:0] <= rx_byte;
                        state <= CHECKSUM_H;
                    end
                    
                    CHECKSUM_H: begin
                        checksum[15:8] <= rx_byte;
                        checksum_valid <= 1'b1;
                        checksum_ok <= (computed_checksum == {rx_byte, checksum[7:0]});
                        state <= IDLE;
                    end
                    
                    default: state <= IDLE;
                endcase
            end
            
            if (packet_end && state != CHECKSUM_H) begin
                state <= IDLE;
                checksum_valid <= 1'b0;
            end
        end
    end
endmodule