//SystemVerilog
module CAN_Interrupt_Controller #(
    parameter DATA_WIDTH = 8
)(
    input clk,
    input rst_n,
    input can_rx,
    output reg can_tx,
    input [DATA_WIDTH-1:0] tx_data,
    input tx_data_valid,
    output reg [DATA_WIDTH-1:0] rx_data,
    output reg tx_irq,
    output reg rx_irq,
    output reg error_irq
);
    reg [2:0] state;
    reg [DATA_WIDTH-1:0] tx_shift;
    reg [3:0] bit_cnt;
    reg rx_active;

    // Added register buffer for bit_cnt to potentially reduce fanout load
    reg [3:0] bit_cnt_buf;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= 0;
            tx_irq <= 0;
            rx_irq <= 0;
            error_irq <= 0;
            bit_cnt <= 0;
            can_tx <= 1'b1;
            tx_shift <= 0;
            rx_data <= 0;
            rx_active <= 0;
            // Reset the buffer register
            bit_cnt_buf <= 0;
        end else begin
            // Update the buffer register with the current bit_cnt value
            // This provides a registered version of bit_cnt that synthesis tools
            // can potentially use to balance fanout or timing paths.
            bit_cnt_buf <= bit_cnt;

            // Original state machine logic remains functionally the same
            case(state)
                0: begin
                    if (can_rx == 1'b0) begin
                        state <= 1;
                        rx_active <= 1;
                        bit_cnt <= 0; // Reset bit counter
                    end
                end
                1: begin
                    rx_data <= {rx_data[DATA_WIDTH-2:0], can_rx};
                    // Original logic using bit_cnt
                    if (bit_cnt == DATA_WIDTH-1) begin
                        rx_irq <= 1;
                        state <= 0;
                        rx_active <= 0;
                    end
                    // Original logic using bit_cnt
                    bit_cnt <= bit_cnt + 1;
                end
                2: begin
                    can_tx <= tx_shift[DATA_WIDTH-1];
                    tx_shift <= {tx_shift[DATA_WIDTH-2:0], 1'b0};
                    // Original logic using bit_cnt
                    if (bit_cnt == DATA_WIDTH-1) begin
                        tx_irq <= 1;
                        state <= 0;
                    end else begin
                        // Original logic using bit_cnt
                        bit_cnt <= bit_cnt + 1;
                    end
                end
                default: begin
                    state <= 0; // Return to idle state
                end
            endcase

            // tx_data_valid logic
            if (tx_data_valid) begin
                tx_shift <= tx_data;
                state <= 2;
                bit_cnt <= 0; // Initialize bit counter
                tx_irq <= 0; // Clear interrupt flag
            end
        end
    end

endmodule