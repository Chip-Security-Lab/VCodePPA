//SystemVerilog
// Half Adder Module
// Adds two 1-bit inputs, produces a sum and a carry-out
module half_adder (
  input wire a,
  input wire b,
  output wire sum,
  output wire carry
);

  assign sum = a ^ b;
  assign carry = a & b;

endmodule

// Full Adder Module
// Adds three 1-bit inputs (a, b, carry-in), produces a sum and a carry-out
module full_adder (
  input wire a,
  input wire b,
  input wire cin,
  output wire sum,
  output wire cout
);

  assign sum = a ^ b ^ cin;
  assign cout = (a & b) | (cin & (a ^ b));

endmodule

// Top-level 2-bit Adder with Structured Data Path
// Instantiates half-adder and full-adder submodules for ripple-carry addition
// Data flow is made explicit through signal naming
module structured_2bit_adder (
  input wire [1:0] data_a,
  input wire [1:0] data_b,
  output wire [2:0] summation
);

  // Internal signals representing the sum and carry output of each stage
  wire stage0_sum;
  wire stage0_carry_out; // Carry-out from LSB stage (Bit 0)

  wire stage1_sum;
  wire stage1_carry_out; // Carry-out from MSB stage (Bit 1)

  // Stage 0 (LSB): Half Adder
  // Adds data_a[0] and data_b[0]
  half_adder u_stage0_adder (
    .a     (data_a[0]),
    .b     (data_b[0]),
    .sum   (stage0_sum),       // Sum for bit 0
    .carry (stage0_carry_out)  // Carry generated by bit 0
  );

  // Stage 1 (MSB): Full Adder
  // Adds data_a[1], data_b[1], and the carry from Stage 0
  full_adder u_stage1_adder (
    .a    (data_a[1]),
    .b    (data_b[1]),
    .cin  (stage0_carry_out), // Carry-in for bit 1 comes from bit 0's carry-out
    .sum  (stage1_sum),       // Sum for bit 1
    .cout (stage1_carry_out)  // Carry generated by bit 1 (final carry-out)
  );

  // Assign the stage outputs to the final summation output array
  // summation[0] is the sum from Stage 0 (LSB)
  // summation[1] is the sum from Stage 1 (MSB)
  // summation[2] is the carry-out from Stage 1 (Most Significant Bit of result)
  assign summation[0] = stage0_sum;
  assign summation[1] = stage1_sum;
  assign summation[2] = stage1_carry_out;

endmodule