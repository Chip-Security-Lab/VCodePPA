//SystemVerilog
module sync_quadrupole_ram_two_write #(
    parameter DATA_WIDTH = 8,
    parameter ADDR_WIDTH = 8
)(
    input wire clk,
    input wire rst,
    input wire we_a, we_b, we_c, we_d,
    input wire [ADDR_WIDTH-1:0] addr_a, addr_b, addr_c, addr_d,
    input wire [DATA_WIDTH-1:0] din_a, din_b, din_c, din_d,
    output reg [DATA_WIDTH-1:0] dout_a, dout_b, dout_c, dout_d
);

    // RAM memory
    reg [DATA_WIDTH-1:0] ram [(2**ADDR_WIDTH)-1:0];
    
    // Pipeline stage 1 - Address and write enable registers
    reg [ADDR_WIDTH-1:0] addr_a_stage1, addr_b_stage1, addr_c_stage1, addr_d_stage1;
    reg [DATA_WIDTH-1:0] din_a_stage1, din_b_stage1, din_c_stage1, din_d_stage1;
    reg we_a_stage1, we_b_stage1, we_c_stage1, we_d_stage1;
    
    // Pipeline stage 2 - RAM read data registers
    reg [DATA_WIDTH-1:0] ram_data_a_stage2, ram_data_b_stage2, ram_data_c_stage2, ram_data_d_stage2;
    reg [ADDR_WIDTH-1:0] addr_a_stage2, addr_b_stage2, addr_c_stage2, addr_d_stage2;
    reg [DATA_WIDTH-1:0] din_a_stage2, din_b_stage2, din_c_stage2, din_d_stage2;
    reg we_a_stage2, we_b_stage2, we_c_stage2, we_d_stage2;
    
    // Pipeline stage 3 - Subtraction result registers
    reg [DATA_WIDTH-1:0] sub_result_a_stage3, sub_result_b_stage3, sub_result_c_stage3, sub_result_d_stage3;
    reg [ADDR_WIDTH-1:0] addr_a_stage3, addr_b_stage3, addr_c_stage3, addr_d_stage3;
    reg we_a_stage3, we_b_stage3, we_c_stage3, we_d_stage3;

    // Stage 1: Register inputs
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            addr_a_stage1 <= 0;
            addr_b_stage1 <= 0;
            addr_c_stage1 <= 0;
            addr_d_stage1 <= 0;
            din_a_stage1 <= 0;
            din_b_stage1 <= 0;
            din_c_stage1 <= 0;
            din_d_stage1 <= 0;
            we_a_stage1 <= 0;
            we_b_stage1 <= 0;
            we_c_stage1 <= 0;
            we_d_stage1 <= 0;
        end else begin
            addr_a_stage1 <= addr_a;
            addr_b_stage1 <= addr_b;
            addr_c_stage1 <= addr_c;
            addr_d_stage1 <= addr_d;
            din_a_stage1 <= din_a;
            din_b_stage1 <= din_b;
            din_c_stage1 <= din_c;
            din_d_stage1 <= din_d;
            we_a_stage1 <= we_a;
            we_b_stage1 <= we_b;
            we_c_stage1 <= we_c;
            we_d_stage1 <= we_d;
        end
    end

    // Stage 2: RAM read
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            ram_data_a_stage2 <= 0;
            ram_data_b_stage2 <= 0;
            ram_data_c_stage2 <= 0;
            ram_data_d_stage2 <= 0;
            addr_a_stage2 <= 0;
            addr_b_stage2 <= 0;
            addr_c_stage2 <= 0;
            addr_d_stage2 <= 0;
            din_a_stage2 <= 0;
            din_b_stage2 <= 0;
            din_c_stage2 <= 0;
            din_d_stage2 <= 0;
            we_a_stage2 <= 0;
            we_b_stage2 <= 0;
            we_c_stage2 <= 0;
            we_d_stage2 <= 0;
        end else begin
            ram_data_a_stage2 <= ram[addr_a_stage1];
            ram_data_b_stage2 <= ram[addr_b_stage1];
            ram_data_c_stage2 <= ram[addr_c_stage1];
            ram_data_d_stage2 <= ram[addr_d_stage1];
            addr_a_stage2 <= addr_a_stage1;
            addr_b_stage2 <= addr_b_stage1;
            addr_c_stage2 <= addr_c_stage1;
            addr_d_stage2 <= addr_d_stage1;
            din_a_stage2 <= din_a_stage1;
            din_b_stage2 <= din_b_stage1;
            din_c_stage2 <= din_c_stage1;
            din_d_stage2 <= din_d_stage1;
            we_a_stage2 <= we_a_stage1;
            we_b_stage2 <= we_b_stage1;
            we_c_stage2 <= we_c_stage1;
            we_d_stage2 <= we_d_stage1;
        end
    end

    // Stage 3: Subtraction
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            sub_result_a_stage3 <= 0;
            sub_result_b_stage3 <= 0;
            sub_result_c_stage3 <= 0;
            sub_result_d_stage3 <= 0;
            addr_a_stage3 <= 0;
            addr_b_stage3 <= 0;
            addr_c_stage3 <= 0;
            addr_d_stage3 <= 0;
            we_a_stage3 <= 0;
            we_b_stage3 <= 0;
            we_c_stage3 <= 0;
            we_d_stage3 <= 0;
        end else begin
            sub_result_a_stage3 <= ram_data_a_stage2 - din_a_stage2;
            sub_result_b_stage3 <= ram_data_b_stage2 - din_b_stage2;
            sub_result_c_stage3 <= ram_data_c_stage2 - din_c_stage2;
            sub_result_d_stage3 <= ram_data_d_stage2 - din_d_stage2;
            addr_a_stage3 <= addr_a_stage2;
            addr_b_stage3 <= addr_b_stage2;
            addr_c_stage3 <= addr_c_stage2;
            addr_d_stage3 <= addr_d_stage2;
            we_a_stage3 <= we_a_stage2;
            we_b_stage3 <= we_b_stage2;
            we_c_stage3 <= we_c_stage2;
            we_d_stage3 <= we_d_stage2;
        end
    end

    // Stage 4: Write back and output
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            dout_a <= 0;
            dout_b <= 0;
            dout_c <= 0;
            dout_d <= 0;
        end else begin
            if (we_a_stage3) ram[addr_a_stage3] <= sub_result_a_stage3;
            if (we_b_stage3) ram[addr_b_stage3] <= sub_result_b_stage3;
            if (we_c_stage3) ram[addr_c_stage3] <= sub_result_c_stage3;
            if (we_d_stage3) ram[addr_d_stage3] <= sub_result_d_stage3;

            dout_a <= ram_data_a_stage2;
            dout_b <= ram_data_b_stage2;
            dout_c <= ram_data_c_stage2;
            dout_d <= ram_data_d_stage2;
        end
    end

endmodule