module add1(input[3:0]x,y, output[4:0]s); 
  assign s = x + y; //4-bit inputs, 5-bit sum
endmodule