//SystemVerilog
module sync_dual_port_ram #(
    parameter DATA_WIDTH = 8,
    parameter ADDR_WIDTH = 8
)(
    input wire clk,
    input wire rst,
    input wire we_a, we_b,
    input wire [ADDR_WIDTH-1:0] addr_a, addr_b,
    input wire [DATA_WIDTH-1:0] din_a, din_b,
    output reg [DATA_WIDTH-1:0] dout_a, dout_b
);

    reg [DATA_WIDTH-1:0] ram [(2**ADDR_WIDTH)-1:0];
    
    // Stage 1: Input registers
    reg [ADDR_WIDTH-1:0] addr_a_stage1, addr_b_stage1;
    reg we_a_stage1, we_b_stage1;
    reg [DATA_WIDTH-1:0] din_a_stage1, din_b_stage1;
    
    // Stage 2: RAM access
    reg [DATA_WIDTH-1:0] ram_data_a_stage2, ram_data_b_stage2;
    reg [ADDR_WIDTH-1:0] addr_a_stage2, addr_b_stage2;
    reg we_a_stage2, we_b_stage2;
    reg [DATA_WIDTH-1:0] din_a_stage2, din_b_stage2;
    
    // Stage 3: Output registers
    reg [DATA_WIDTH-1:0] ram_data_a_stage3, ram_data_b_stage3;

    // Stage 1: Input pipeline
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            addr_a_stage1 <= 0;
            addr_b_stage1 <= 0;
            we_a_stage1 <= 0;
            we_b_stage1 <= 0;
            din_a_stage1 <= 0;
            din_b_stage1 <= 0;
        end else begin
            addr_a_stage1 <= addr_a;
            addr_b_stage1 <= addr_b;
            we_a_stage1 <= we_a;
            we_b_stage1 <= we_b;
            din_a_stage1 <= din_a;
            din_b_stage1 <= din_b;
        end
    end

    // Stage 2: RAM access pipeline
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            ram_data_a_stage2 <= 0;
            ram_data_b_stage2 <= 0;
            addr_a_stage2 <= 0;
            addr_b_stage2 <= 0;
            we_a_stage2 <= 0;
            we_b_stage2 <= 0;
            din_a_stage2 <= 0;
            din_b_stage2 <= 0;
        end else begin
            addr_a_stage2 <= addr_a_stage1;
            addr_b_stage2 <= addr_b_stage1;
            we_a_stage2 <= we_a_stage1;
            we_b_stage2 <= we_b_stage1;
            din_a_stage2 <= din_a_stage1;
            din_b_stage2 <= din_b_stage1;
            
            if (we_a_stage1) ram[addr_a_stage1] <= din_a_stage1;
            if (we_b_stage1) ram[addr_b_stage1] <= din_b_stage1;
            
            ram_data_a_stage2 <= ram[addr_a_stage1];
            ram_data_b_stage2 <= ram[addr_b_stage1];
        end
    end

    // Stage 3: Output pipeline
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            ram_data_a_stage3 <= 0;
            ram_data_b_stage3 <= 0;
        end else begin
            ram_data_a_stage3 <= ram_data_a_stage2;
            ram_data_b_stage3 <= ram_data_b_stage2;
        end
    end

    // Output assignment
    assign dout_a = ram_data_a_stage3;
    assign dout_b = ram_data_b_stage3;

endmodule