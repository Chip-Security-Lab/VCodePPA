//SystemVerilog
module adder_8bit_cla (
  input [7:0] a,
  input [7:0] b,
  input       cin,
  output [7:0] sum,
  output      cout
);

  wire [7:0] p; // propagate: a_i ^ b_i
  wire [7:0] g; // generate: a_i & b_i

  assign p = a ^ b;
  assign g = a & b;

  // Internal carries (c[0] is cin, c[i] is carry into bit i for i=1..7)
  // c[8] is the final carry out (cout)
  wire [8:0] c;

  // Input carry
  assign c[0] = cin;

  // Full 8-bit Carry Lookahead Logic (fully expanded)
  // c[i+1] = g[i] | (p[i] & g[i-1]) | (p[i] & p[i-1] & g[i-2]) | ... | (p[i] & ... & p[0] & c[0])
  assign c[1] = g[0] | (p[0] & c[0]);
  assign c[2] = g[1] | (p[1] & g[0]) | (p[1] & p[0] & c[0]);
  assign c[3] = g[2] | (p[2] & g[1]) | (p[2] & p[1] & g[0]) | (p[2] & p[1] & p[0] & c[0]);
  assign c[4] = g[3] | (p[3] & g[2]) | (p[3] & p[2] & g[1]) | (p[3] & p[2] & p[1] & g[0]) | (p[3] & p[2] & p[1] & p[0] & c[0]);
  assign c[5] = g[4] | (p[4] & g[3]) | (p[4] & p[3] & g[2]) | (p[4] & p[3] & p[2] & g[1]) | (p[4] & p[3] & p[2] & p[1] & g[0]) | (p[4] & p[3] & p[2] & p[1] & p[0] & c[0]);
  assign c[6] = g[5] | (p[5] & g[4]) | (p[5] & p[4] & g[3]) | (p[5] & p[4] & p[3] & g[2]) | (p[5] & p[4] & p[3] & p[2] & g[1]) | (p[5] & p[4] & p[3] & p[2] & p[1] & g[0]) | (p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & c[0]);
  assign c[7] = g[6] | (p[6] & g[5]) | (p[6] & p[5] & g[4]) | (p[6] & p[5] & p[4] & g[3]) | (p[6] & p[5] & p[4] & p[3] & g[2]) | (p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]) | (p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & c[0]);
  assign c[8] = g[7] | (p[7] & g[6]) | (p[7] & p[6] & g[5]) | (p[7] & p[6] & p[5] & g[4]) | (p[7] & p[6] & p[5] & p[4] & g[3]) | (p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]) | (p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & c[0]);

  // Sum bits calculation
  // sum[i] = p[i] ^ c[i]
  assign sum[0] = p[0] ^ c[0];
  assign sum[1] = p[1] ^ c[1];
  assign sum[2] = p[2] ^ c[2];
  assign sum[3] = p[3] ^ c[3];
  assign sum[4] = p[4] ^ c[4];
  assign sum[5] = p[5] ^ c[5];
  assign sum[6] = p[6] ^ c[6];
  assign sum[7] = p[7] ^ c[7];

  // Final carry out
  assign cout = c[8];

endmodule