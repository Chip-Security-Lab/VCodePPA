module xor_base(input a, b, output y);
    assign y = a ^ b;
endmodule