module TriStateNOT(
    input oe,  // Output enable
    input [3:0] in,
    output [3:0] out
);
    assign out = oe ? ~in : 4'bzzzz;
endmodule
