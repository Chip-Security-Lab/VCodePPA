module adder_2 (input x, y, output z);
  assign z = x + y;
endmodule