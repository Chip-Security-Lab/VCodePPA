module AND_Basic(
    input a, b,
    output y
);
    assign y = a & b; // 基础两输入与门
endmodule
